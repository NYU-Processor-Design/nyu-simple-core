module Core;


endmodule
